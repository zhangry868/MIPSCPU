module InstruMemory 
#(parameter DATA_WIDTH = 32, parameter ADDR_WIDTH = 32)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input [3:0] we, 
	input clk,
	output [(DATA_WIDTH-1):0] q
);

	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] ram[2**(ADDR_WIDTH - 22) - 1:0];

	// Variable to hold the registered read address
	reg [ADDR_WIDTH-1:0] addr_reg;
	
initial
begin
/*
ram[0] = 32'b000000_00010_00011_00011_00000_100000;
ram[1] = 32'b000000_00010_00011_00011_00000_100000;//2# + 3# ->3#
ram[2] = 32'b000000_00010_00001_00010_00000_100010;//2# - 1#
ram[3] = {16'b000001_00010_00010,16'hfffd};//begz 2# > 0
ram[4] = {16'b000001_00011_00011,16'hffff};//begz 3# > 0
*/
//1# 1
//2# 2
//Add Sub

//--------------------------------------------Test1-------------------------------------------

ram[0] = 32'b000000_01001_01010_00011_00000_100000;//3# 3 
ram[1] = 32'b000000_01001_01100_00100_00000_100010;//9# - 12#
ram[2] = 32'b000000_11111_00100_00101_00000_100010;//31# - 4# ->5# Overflow
ram[3] = 32'b000000_00101_00001_00011_00000_100000;//5# + 1# ->5#
//5# 6

ram[4] = 32'b000000_00100_00001_00101_00000_100011;//subu 4# - 1# ->5# 5#ffffffe
ram[5] = 32'b000000_00010_00101_00101_00000_000111;//SRAV 5# >> (2#:2)
ram[6] = 32'b000000_00010_01001_00101_00010_000010;//ROTR 9# >> (Shamat)->5#
ram[7] = 32'b000000_01010_01001_00101_00000_101011;//sltu 10# - 9# -> 5#
//???????5# fffffff
ram[8] = {16'b001000_00101_00101,16'h789a};//addi 5# I ->5#
ram[9] = {16'b001000_11111_00101,16'h7abc};//addi 31# I ->5#  
ram[10] = {16'b001001_11111_00101,16'h7abc};//addiu 31# I ->5#  
ram[11] = {16'b001001_00101_00101,16'h789a};//addiu 5# I ->5#

ram[12] = {16'b001111_00000_00101,16'h789a};//lui lui I ->5#
ram[13] = {16'b001110_11111_00101,16'habcd};//xori xori I 31# -> 5#

ram[14] = 32'b011100_01011_00010_00101_00000_100001;//clo 11# ->5#
ram[15] = 32'b011100_01010_00010_00101_00000_100000;//clz 10# ->5#
ram[16] = {16'b001010_00101_00101,16'habcd};//slti  5# < I ->5#
ram[17] = 32'b011111_00000_01101_00110_10000_100000;//seb 8# -> 6#
ram[18] = {16'b101011_00000_01001,16'd512};//sw
ram[19] = {16'b101010_00000_11111,16'd256};//swl
ram[20] = {16'b100011_00000_00011,16'd512};//lw
ram[21] = {16'b100010_00000_00011,16'd513};//lwl
ram[22] = {16'b100010_00000_00011,16'd514};//lwl
ram[23] = {16'b100010_00000_00011,16'd515};//lwl
ram[24] = {16'b100110_00000_00011,16'd513};//lwr
ram[25] = {16'b100110_00000_00011,16'd514};//lwr
ram[26] = {16'b100110_00000_00011,16'd515};//lwr
ram[27] = 32'b000000_01001_00011_00011_00000_100000;//3# 3 
//ram[8'b10000000] = 32'h7fffffff;
ram[28] = {16'b101010_00000_11111,16'd513};//swl
ram[29] = {16'b101010_00000_11111,16'd514};//swl
ram[30] = {16'b101010_00000_11111,16'd515};//swl
ram[31] = {16'b101110_00000_11111,16'd513};//swr
ram[32] = {16'b101110_00000_11111,16'd514};//swr
ram[33] = {16'b101110_00000_11111,16'd515};//swr
ram[34] = {16'b000001_00001_10001,16'h0006};//begzal 1# > 0
//ram[19] = {16'b000001_00001_00001,16'h0010};//begz 1# > 0
ram[35] = {6'b000010,2'b0,24'h0};//J
ram[41] = {16'b000001_11110_00001,16'h0001};//begz 30# < 0

ram[42] = {6'b000010,2'b0,24'h0};//J


//-------------------------Test2--------------------------------------------------------------
//ram[0] = {16'b101011_00000_01001,16'd512};//sw
//ram[1] = {16'b100011_00000_01110,16'd512};//lw
//ram[2] = 32'b000000_01110_00001_00001_00000_100000;
/*
ram[0] = 32'b0;
ram[1] = 32'b0;
ram[2] = 32'b0;
ram[3] = 32'b0;
ram[4] = {16'b101011_00000_01001,16'd512};//sw
ram[5] = {16'b101010_00000_11111,16'd256};//swl
ram[6] = {16'b100011_00000_00011,16'd512};//lw
ram[7] = {16'b100010_00000_00011,16'd513};//lwl
ram[8] = {16'b100010_00000_00011,16'd514};//lwl
ram[9] = {16'b100010_00000_00011,16'd515};//lwl
ram[10] = {16'b100110_00000_00011,16'd513};//lwr
ram[11] = {16'b100110_00000_00011,16'd514};//lwr
ram[12] = {16'b100110_00000_00011,16'd515};//lwr
//ram[8'b10000000] = 32'h7fffffff;
ram[13] = {16'b101010_00000_11111,16'd513};//swl
ram[14] = {16'b101010_00000_11111,16'd514};//swl
ram[15] = {16'b101010_00000_11111,16'd515};//swl
ram[16] = {16'b101110_00000_11111,16'd513};//swr
ram[17] = {16'b101110_00000_11111,16'd514};//swr
ram[18] = {16'b101110_00000_11111,16'd515};//swr
*/

//----------------------------Test3----------------------------------------------------------
/*ram[0] = {16'b000001_11111_10001,16'd10};//bgezal
//ram[1] = {16'b000001_11111_00001,16'hffff};//begz 3# > 0
ram[2] = {16'b000001_11111_00001,16'hffff};//begz 3# > 0
ram[11] = {16'b000001_11111_00001,16'hffff};//begz 3# > 0*/
//----------------------------Test4----------------------------------------------------------
/*ram[0] = 32'b000000_00010_00011_00011_00000_100000;//2# + 3# ->3#
ram[1] = 32'b000000_00010_00001_00010_00000_100010;//2# - 1#
ram[2] = {16'b000001_00010_00001,16'hfffd};//begz 2# > 0
ram[3] = {16'b000001_00011_00001,16'hffff};//begz 3# > 0
*/
//----------------------------Test5----------------------------------------------------------
/*
ram[0] = 32'h00644020;        //1 - add r8 = r3 + r4 不溢出
ram[1] = 32'h00654020;        //1 - add r8 = r3 + r5 溢出
ram[2] = 32'h20670000;        //2 -addi r7  = r3 + 0000 不溢出
ram[3] = 32'h2027fffe;        //2 -addi r7  = r1 + fffe 溢出
ram[4] = 32'h2426fffe;        //3 -addiu r6 = r1 + fffe 溢出但不判断不溢出
ram[5] = 32'h00694022;        //4 -sub   r8 = r3 - r9  不溢出
ram[6] = 32'h006a6022;        //4 -sub   r12 = r3 - r10  溢出
ram[7] = 32'h006a6023;        //5 -subu  r12 = r3 - r10  溢出但不溢出
ram[8] = 32'h7c0b6420;        //6 -seb   r12 = r11 第八位符号扩展
ram[9] = 32'h3c0d1234;        //7 -lui   r13 = im 低位存入高位 
ram[10] = 32'h38670000;       //8 -xori  r7 = r3 nor im
ram[11] = 32'h70804021;       //9 -clo   r8 = r4 前导1 *rd_in
ram[12] = 32'h70604020;       //10 -clz  r8 = r3 前导0 *rd
ram[13] = 32'h004b4007;       //11 -srav r8 = r11 右移移动 r2位

ram[14] = 32'h002b40c2;       //12 -rotr r8 = r11 右移移动 shamt =3 位
ram[15] = 32'h0043402b;       //13 -sltu r2 r3 比较大小 结果存入r8  
ram[16] = 32'h28480000;       //14 -slti r2 im 比较大小 结果存入r8
ram[17] = 32'h28480fff;       //14 -slti r2 im 比较大小 结果存入r8
ram[18] = 32'h08000020;       //15 -j 跳转到 32 
ram[32] = 32'h04400004;       //16 -bgezal  r2 大于等于0 则跳转 offset<<2  save r31 
	
ram[36] = 32'h880800e1;       //18 -lwl r0+im(56)代表的寄存器值移位(8)后存入r8
ram[37] = 32'h8c0800e0;       //19 -lw  r0+im(56)代表的寄存器值移位(0)后存入r8	
ram[38] = 32'hac0400e0;       //20 -sw  r0+im(56)代表的内存存入R4移位(0)后的值
ram[39] = 32'hb80400e1;       //21 -swr r0+im(56)代表的内存存入R4移位(8)后的值
	
//process-1
ram[40] = 32'h8c0200e4;       //19 -lw  r0+im(57)代表的寄存器值移位(0)后存入r2  
											//r2计数器置为-5
ram[41] = 32'h00004020;       //1 - add r8 = r0 + r0     r8清零	
ram[42] = 32'h20420001;       //2 -addi r2 = r2 + 0001   计数器+1  
ram[43] = 32'h04400004;       //16 -bgezal  r2 大于等于0 则跳转 offset<<2  save r31 
											//r2>=0后跳出循环
ram[44] = 32'hac0200e0;       //20 -sw  r0+im(56)代表的内存存入R2移位(0)后的值
ram[45] = 32'h0800002a;       //15 -j 跳转到 42 

ram[56] = 32'h0f0f0f0f;
ram[57] = 32'hfffffffa;	
*/
/*
ram[0] = 32'b001000_00000_00111_0000000000000100;  //addi r0 im(4) -> r7
ram[1] = 32'b000000_00000_00111_0100000000100010;  //sub  r0 r7 -> r8
ram[2] = 32'b001000_01000_01000_0000000000000001;  //addi r8 im(1) -> r8

ram[3] = 32'b000000_00010_00001_0101000000100010;  //sub  r2 r1 -> r10
ram[4] = 32'b000001_01010_00001_0000000000000011; //bgez r10 -> 3
ram[5] = 32'b000000_00000_00001_0100100000100111; //nor r0 r1 -> r9
ram[6] = 32'b000000_00000_00010_0000100000100111; //nor r0 r2 -> r1
ram[7] = 32'b000000_00000_01001_0001000000100111; //nor r0 r9 -> r2

ram[8] = 32'b000000_00011_00010_0101000000100010;  //sub  r3 r2 -> r10
ram[9] = 32'b000001_01010_00001_0000000000000011; //bgez r10 -> 3
ram[10] = 32'b000000_00000_00010_0100100000100111; //nor r0 r2 -> r9
ram[11] = 32'b000000_00000_00011_0001000000100111; //nor r0 r3 -> r2
ram[12] = 32'b000000_00000_01001_0001100000100111; //nor r0 r9 -> r3

ram[13] = 32'b000000_00100_00011_0101000000100010;  //sub  r4 r3 -> r10
ram[14] = 32'b000001_01010_00001_0000000000000011; //bgez r10 -> 3
ram[15] = 32'b000000_00000_00011_0100100000100111; //nor r0 r3 -> r9
ram[16] = 32'b000000_00000_00100_0001100000100111; //nor r0 r4 -> r3
ram[17] = 32'b000000_00000_01001_0010000000100111; //nor r0 r9 -> r4

ram[18] = 32'b000000_00101_00100_0101000000100010;  //sub  r5 r4 -> r10
ram[19] = 32'b000001_01010_00001_0000000000000011; //bgez r10 -> 3
ram[20] = 32'b000000_00000_00100_0100100000100111; //nor r0 r4 -> r9
ram[21] = 32'b000000_00000_00101_0010000000100111; //nor r0 r5 -> r4
ram[22] = 32'b000000_00000_01001_0010100000100111; //nor r0 r9 -> r5

ram[23] = 32'b000001_01000_00001_0000000000000001; //bgez r8 -> 1
ram[24] = 32'b000010_00000_00000_0000000000000010; //j    jump to 2
*/
end
	
	always @ (negedge clk)
	begin
		// Write
		if (we[0] == 1'b1)
			ram[addr[9:2]][7:0] <= data[7:0];
		if (we[1] == 1'b1)
			ram[addr[9:2]][15:8] <= data[15:8];
		if (we[2] == 1'b1)
			ram[addr[9:2]][23:16] <= data[23:16];
		if (we[3] == 1'b1)
			ram[addr[9:2]][31:24] <= data[31:24];
		//addr_reg <= addr;
	end
	
	// Continuous assignment implies read returns NEW data.
	// This is the natural behavior of the TriMatrix memory
	// blocks in Single Port mode.  
	assign q = ram[addr[9:2]];

endmodule
