library verilog;
use verilog.vl_types.all;
entity ID_EX_Seg is
    port(
        Clk             : in     vl_logic;
        stall           : in     vl_logic;
        flush           : in     vl_logic;
        PC_Add          : in     vl_logic_vector(31 downto 0);
        OverflowEn      : in     vl_logic;
        condition       : in     vl_logic_vector(2 downto 0);
        Branch          : in     vl_logic;
        PC_write        : in     vl_logic_vector(2 downto 0);
        Mem_Byte_Write  : in     vl_logic_vector(3 downto 0);
        Rd_Write_Byte_en: in     vl_logic_vector(3 downto 0);
        MemWBSrc        : in     vl_logic;
        Jump            : in     vl_logic;
        ALUShiftSrc     : in     vl_logic;
        MemDataSrc      : in     vl_logic_vector(2 downto 0);
        ALUSrcA         : in     vl_logic;
        ALUSrcB         : in     vl_logic;
        ALUOp           : in     vl_logic_vector(3 downto 0);
        RegDst          : in     vl_logic_vector(1 downto 0);
        ShiftAmountSrc  : in     vl_logic;
        ShiftOp         : in     vl_logic_vector(1 downto 0);
        OperandA        : in     vl_logic_vector(31 downto 0);
        OperandB        : in     vl_logic_vector(31 downto 0);
        Rs              : in     vl_logic_vector(4 downto 0);
        Rt              : in     vl_logic_vector(4 downto 0);
        Rd              : in     vl_logic_vector(4 downto 0);
        Immediate32     : in     vl_logic_vector(31 downto 0);
        Shamt           : in     vl_logic_vector(4 downto 0);
        BranchSel       : in     vl_logic;
        RtRead          : in     vl_logic_vector(1 downto 0);
        PC_Add_out      : out    vl_logic_vector(31 downto 0);
        OverflowEn_out  : out    vl_logic;
        condition_out   : out    vl_logic_vector(2 downto 0);
        Branch_out      : out    vl_logic;
        PC_write_out    : out    vl_logic_vector(2 downto 0);
        Mem_Byte_Write_out: out    vl_logic_vector(3 downto 0);
        Rd_Write_Byte_en_out: out    vl_logic_vector(3 downto 0);
        MemWBSrc_out    : out    vl_logic;
        Jump_out        : out    vl_logic;
        ALUShiftSrc_out : out    vl_logic;
        MemDataSrc_out  : out    vl_logic_vector(2 downto 0);
        ALUSrcA_out     : out    vl_logic;
        ALUSrcB_out     : out    vl_logic;
        ALUOp_out       : out    vl_logic_vector(3 downto 0);
        RegDst_out      : out    vl_logic_vector(1 downto 0);
        ShiftAmountSrc_out: out    vl_logic;
        ShiftOp_out     : out    vl_logic_vector(1 downto 0);
        OperandA_out    : out    vl_logic_vector(31 downto 0);
        OperandB_out    : out    vl_logic_vector(31 downto 0);
        Rs_out          : out    vl_logic_vector(4 downto 0);
        Rt_out          : out    vl_logic_vector(4 downto 0);
        Rd_out          : out    vl_logic_vector(4 downto 0);
        Immediate32_out : out    vl_logic_vector(31 downto 0);
        Shamt_out       : out    vl_logic_vector(4 downto 0);
        BranchSel_out   : out    vl_logic;
        RtRead_out      : out    vl_logic_vector(1 downto 0)
    );
end ID_EX_Seg;
