library verilog;
use verilog.vl_types.all;
entity pipeline_vlg_tst is
end pipeline_vlg_tst;
